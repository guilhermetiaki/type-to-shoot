library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity ger_palavras is
	port ( KEY 	:		in	STD_LOGIC_VECTOR (3 downto 0);		--	Pushbutton[3:0]
			 PS2_DAT 	:		inout	STD_LOGIC;	--	PS2 Data
		    PS2_CLK		:		inout	STD_LOGIC;		--	PS2 Clock
			 CLOCK_24	: 	in	STD_LOGIC_VECTOR (1 downto 0);	--	24 MHz
	       clk : in std_logic;
			 init_line: out integer range 0 to 95;

			 init_col: out INTEGER range 0 to 56;

			 reset : buffer STD_LOGIC;

			 mapaLetras : buffer STD_LOGIC_VECTOR (0 to 299);
			
			 LEDG 	:		out	STD_LOGIC_VECTOR (7 downto 0);
			 LEDR 	:		out	STD_LOGIC_VECTOR (9 downto 0)
			);
end ger_palavras;

architecture comportamento of ger_palavras is

	component kbdex_ctrl
		generic(
			clkfreq : integer
		);
		port(
			ps2_data	:	inout	std_logic;
			ps2_clk		:	inout	std_logic;
			clk				:	in 	std_logic;
			en				:	in 	std_logic;
			resetn		:	in 	std_logic;
			lights		: in	std_logic_vector(2 downto 0); -- lights(Caps, Nun, Scroll)		
			key_on		:	out	std_logic_vector(2 downto 0);
			key_code	:	out	std_logic_vector(47 downto 0)
		);
	end component;
	
	component mapeador
		port(
			letra : in std_logic_vector(4 downto 0);
			mapa : out std_logic_vector(0 to 24)
		);
	end component;


	SIGNAL enable: STD_LOGIC; -- sinal que avisa pra pegar o contador de rangom gen

	SIGNAL slow_clock: STD_LOGIC;
	
	SIGNAL start_screen: STD_LOGIC;
	
	SIGNAL CLOCK_DIV : INTEGER := 5000000;

	SIGNAL palavras : STD_LOGIC_VECTOR (0 to 2999);
	signal codigoLetras : STD_LOGIC_VECTOR (0 to 1919);
	
	signal index: integer range 0 to 56;
	
	signal index2: integer range 0 to 9;

	
	signal letrasComidas: integer range 0 to 12;
	signal palavrasComidas: integer range 0 to 9;
	
	signal arrh :std_LOGIC;
	
	signal keys_on :std_LOGIC;
	
	signal palavra_digitada: STD_LOGIC;
	
	signal line: integer range 0 to 95;

	signal key_on	: std_logic_vector( 2 downto 0);
	signal key0 : std_logic_vector(15 downto 0);
	
begin
	palavras <= "100011000111111100011000111110100011111010000100001111010001111101000010000111111000011110100001111101110100011111110001100011111110001111111001010001111111000011110100001111111110100011000110001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101000111110100011111011111100011111110010100011111100100001000010011111011101000010011100010111010001100011111110001100011111100100001000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000010000100001111111111001000010000100111111111100100001000010000100111111000011110100001111111111100011111110010100010111010001111111000110001100001000010000100001111110000100001000010000111111000111011011100010001100000000000000000000000000000000000000000000000000000000000000000000000000000111110010000100001001111110001110011010110011100011000110001010100101000100011101000111111100011000110000100001000010000111111111100100001000010011111111101000110001100011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101000110001100010111011110100011111010001111100001100001000011000101110111111000011110100001111101110100011000010001011101111100100001000010000100111110010000100001001111101110100011000110001011101000111001101011001110001000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111100101000111111100001111010000111111000111011101011000110001111111000011110100001111110001110111010110001100011111010001111101000111110111111000011110100001111111111100011111110010100011111110000111101000011111111101000110001100011111000000000000000000000000000000000000000000000000000111101000110001100011111011111100001111010000111111000010000100001000011111111110010000100001001111110001100010101001010001001111110000111101000011111111111000111111100101000111111100001111010000111111111010001100011000111110000000000000000000000000000000000000000000000000000000000000000000000000000111110010000100001000010011111100011111110010100010111010001111111000110001100011100110101100111000101111100000111000001111101000010000100001000011111011101000111111100011000111111001000010000100001001111100100001000010011111011101000110001100010111010001110011010110011100010000000000000000000000000011101000110001100010111011110100011111010000100001111100100001000010011111100011100110101100111000111111001000010000100111110111010001100011000101110100011100110101100111000101111100000111000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000110001100010111010001110011010110011100011111010001100011000111110111111000011110100001111111111100011111110010100010111110000011100000111110111110010000100001000010001110100011111110001100011000111001101011001110001111101000110001100011111000000000000000000000000000000000000000000000000000";
	
	codigoLetras <= "000000000001110000000000010011010000000001001101000000000010010000000000000111000000000000101101000000000010010000000000001000110000000000000000000000000000000000000000000000000000000000000000000000000011001000000000001011010000000001000011000000000011010000000000001100110000000000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101100000000010000110000000000101100000000000010010000000000001011010000000000011100000000000100101100000000010010110000000000110101000000000000000000000000000000000000000000000000000000000100001100000000001100010000000000101010000000000001110000000000010010110000000001000011000000000010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000001100100000000000111011000000000010010000000000001000010000000000101100000000000100001100000000010001000000000000110001000000000000000000000000000000000000000000000000000000000010110100000000001001000000000000111010000000000010010000000000001110100000000000110010000000000010010000000000001011010000000000100100000000000010001100000000000000000000000000000000000000000010001100000000001001000000000001001011000000000100001100000000001010100000000000100100000000000010110100000000001001000000000000100011000000000000000000000000000000000000000000000000000000000010110000000000001011010000000000011100000000000011000100000000000110110000000001001011000000000001110000000000001011000000000001000011000000000100010000000000001100010000000000000000000000000100010000000000010011010000000001000011000000000011000100000000010000110000000001000100000000000011000100000000000110110000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001100010000000000100011000000000010010000000000001011010000000000011011000000000010110000000000000111000000000000110001000000000010001100000000000000000000000000000000";

	init_line <= line;

	kbd_ctrl : kbdex_ctrl generic map(24000) port map(
		PS2_DAT, PS2_CLK, CLOCK_24(0), key(1), key(0), "000", key_on, key_code(15 downto 0) => key0);
	
	keys_on <= key_on(0) or key_on(1) or key_on(2);
	
	main:
	process (keys_on, palavra_digitada, reset)
	begin
		if(reset = '1') or palavra_digitada = '1' then
			letrasComidas <= 0;
			init_col <= index;
			palavra_digitada <= '0';
		elsif(rising_edge(keys_on)) then
			if(index2 = 0) then
				if(key0 = codigoLetras(letrasComidas*16 to letrasComidas*16 + 15)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 1) then
				if(key0 = codigoLetras(12*16*1+letrasComidas*16 to 12*16*1+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 2) then
				if(key0 = codigoLetras(12*16*2+letrasComidas*16 to 12*16*2+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 3) then
				if(key0 = codigoLetras(12*16*3+letrasComidas*16 to 12*16*3+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 4) then
				if(key0 = codigoLetras(12*16*4+letrasComidas*16 to 12*16*4+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 5) then
				if(key0 = codigoLetras(12*16*5+letrasComidas*16 to 12*16*5+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 6) then
				if(key0 = codigoLetras(12*16*6+letrasComidas*16 to 12*16*6+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 7) then
				if(key0 = codigoLetras(12*16*7+letrasComidas*16 to 12*16*7+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 8) then
				if(key0 = codigoLetras(12*16*8+letrasComidas*16 to 12*16*8+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			elsif(index2 = 9) then
				if(key0 = codigoLetras(12*16*9+letrasComidas*16 to 12*16*9+(letrasComidas+1)*16 - 1)) then
					letrasComidas <= letrasComidas + 1;
				end if;
			end if;
		end if;
		
		
		if letrasComidas = 0 then
			mapaLetras <= palavras(index2*300 to (index2+1)*300 - 1);
		elsif mapaLetras = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" then
			palavra_digitada <= '1';
		else
			mapaLetras(0 to 299) <= palavras(index2*300 to (index2+1)*300 - 1);
			mapaLetras(0 to letrasComidas*25 - 1) <= (OTHERS => '0');
		end if;
	end process;

	move_letra: 
	process (slow_clock)
	begin  -- process conta_coluna;
		if reset = '1' or palavra_digitada = '1' then
			line <= 0;
		elsif slow_clock'event and slow_clock = '1' then  -- rising clock edge
			if line = 90 then               -- conta de 0 a 95 (96 linhas)
				start_screen <= '1';
			else
				line <= line + 2;  
			end if;
		end if;
	
	end process move_letra;
	
	random:
	PROCESS (clk, enable, slow_clock)
		VARIABLE j : INTEGER := 0;
	BEGIN
	
		if(rising_edge(slow_clock)) then
			index <= j;
		end if;

		IF (rising_edge(clk)) THEN
			if j = 56 then      
          j := 0;
			else
          j := j + 1;
			end if;
		END IF;
		
	END PROCESS random;
	
	random2:
	PROCESS (clk, palavra_digitada, reset)
		VARIABLE k : INTEGER := 0;
	BEGIN
		arrh <= palavra_digitada or reset;
		
		if arrh='1' then
			index2 <= k;
		end if;

		IF (rising_edge(clk)) THEN
			if k = 9 then      
          k := 0;
			else
          k := k + 1;
			end if;
		END IF;
		
	END PROCESS random2;
	
	resetatudo:
	process (key(3), key_on(0), line)
	begin
		if key(3) = '0' or line = 90 then
			reset <= '1';
		elsif rising_edge(key_on(0)) then
			reset <= '0';
		end if;
	end process;				  
					  
	clock_divider:
	PROCESS (clk)
		VARIABLE i : INTEGER := 0;
	BEGIN

		IF (rising_edge(clk)) THEN
			IF (i <= CLOCK_DIV/2) THEN
				i := i + 1;
				slow_clock <= '0';
			ELSIF (i < CLOCK_DIV-1) THEN
				i := i + 1;
				slow_clock <= '1';
			ELSE		
				i := 0;
			END IF;	
		END IF;
	END PROCESS;
	
	
end comportamento;