library ieee;
use ieee.std_logic_1164.all;

entity mapeador is
  port (    
    clk27M      : in  std_logic;    
    red, green, blue          : out std_logic_vector(3 downto 0);
    hsync, vsync              : out std_logic;
	 
	PS2_DAT 	:		inout	STD_LOGIC;	--	PS2 Data
	 PS2_CLK		:		inout	STD_LOGIC;		--	PS2 Clock
	 CLOCK_24	: 	in	STD_LOGIC_VECTOR (1 downto 0);	--	24 MHz
	 HEX0 	:		out	STD_LOGIC_VECTOR (6 downto 0);		--	Seven Segment Digit 0
	 KEY 	:		in	STD_LOGIC_VECTOR (3 downto 0);		--	Pushbutton[3:0]
	 
	 
	 LEDG 	:		out	STD_LOGIC_VECTOR (7 downto 0);
	 LEDR 	:		out	STD_LOGIC_VECTOR (9 downto 0)

	 );
end mapeador;

architecture comportamento of mapeador is
  -- Interface com a mem�ria de v�deo do controlador

  signal we : std_logic;                        -- write enable ('1' p/ escrita)
  signal addr : integer range 0 to 12287;       -- endereco mem. vga
  signal pixel : std_logic_vector(2 downto 0);  -- valor de cor do pixel
  signal pixel_bit : std_logic;                 -- um bit do vetor acima

  -- Sinais dos contadores de linhas e colunas utilizados para percorrer
  -- as posi��es da mem�ria de v�deo (pixels) no momento de construir um quadro.
  
  signal line : integer range 0 to 95;  -- linha atual
  signal col : integer range 0 to 127;  -- coluna atual

	signal init_line : integer range 0 to 95;  -- linha atual
	signal init_col : integer range 0 to 127;  -- coluna atual
	
	signal start_screen : STD_LOGIC_VECTOR (0 to 12287) := "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100010111100111110000000111110011100000000011110100010011100011100111110000000000000000000000000000000000000000000000000000010001101101000101000000000000010001000100000001000001000101000101000100010000000000000000000000000000000000000000000000000000000100001110011110011110000000000100010001000000001110011111010001010001000100000000000000000000000000000000000000000000000000000001000001000100000100000000000001000100010000000000010100010100010100010001000000000000000000000000000000000000000000000000000000010000110001000001111100000000010000111000000001111001000100111000111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100111110111110011110011110000000011100100010100010000000100010111110100010000000000000000000000000000000000000000000000000001000101000101000001000001000000000001000101100101101100000001001001000001101100000000000000000000000000000000000000000000000000011110011111011110001110001110000000011111010101001110000000011100011110001110000000000000000000000000000000000000000000000000000100000100100100000000010000010000000100010100110001000000000100100100000001000000000000000000000000000000000000000000000000000001000001000101111101111001111000000001000101000100110000000001000101111100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100111000000000111101111100111001111101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000010000000100010001010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000011100001000111110111110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000000100010001000101001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001110000000011110000100010001010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	
	SIGNAL mapaLetras : STD_LOGIC_VECTOR (0 to 299);
	
	SIGNAL reset : STD_LOGIC;

begin  -- comportamento


  -- Aqui instanciamos o controlador de v�deo, 128 colunas por 96 linhas
  -- (aspect ratio 4:3). Os sinais que iremos utilizar para comunicar
  -- com a mem�ria de v�deo (para alterar o brilho dos pixels) s�o
  -- write_clk (nosso clock), write_enable ('1' quando queremos escrever
  -- o valor de um pixel), write_addr (endere�o do pixel a escrever)
  -- e data_in (valor do brilho do pixel RGB, 1 bit pra cada componente de cor)
  vga_controller: entity work.vgacon port map (
    clk27M       => clk27M,
    rstn         => '1',
    red          => red,
    green        => green,
    blue         => blue,
    hsync        => hsync,
    vsync        => vsync,
    write_clk    => clk27M,
    write_enable => '1',
    write_addr   => addr,
    data_in      => pixel
	 );

  -----------------------------------------------------------------------------
  -- Processos que controlam contadores de linhas e coluna para varrer
  -- todos os endere�os da mem�ria de v�deo, no momento de construir um quadro.
  -----------------------------------------------------------------------------

  -- purpose: Este processo conta o n�mero da coluna atual, quando habilitado
  --          pelo sinal "col_enable".
  -- type   : sequential
  -- inputs : clk27M, col_rstn
  -- outputs: col
  conta_coluna: process (clk27M)
  begin  -- process conta_coluna
    if clk27M'event and clk27M = '1' then  -- rising clock edge
        if col = 127 then               -- conta de 0 a 127 (128 colunas)
          col <= 0;
        else
          col <= col + 1;  
        end if;
    end if;
  end process conta_coluna;
    
  -- purpose: Este processo conta o n�mero da linha atual, quando habilitado
  --          pelo sinal "line_enable".
  -- type   : sequential
  -- inputs : clk27M, line_rstn
  -- outputs: line
  conta_linha: process (clk27M)
  begin  -- process conta_linha
    if clk27M'event and clk27M = '1' then  -- rising clock edge
      -- o contador de linha s� incrementa quando o contador de colunas
      -- chegou ao fim (valor 127)
      if col = 127 then
        if line = 95 then               -- conta de 0 a 95 (96 linhas)
          line <= 0;
        else
          line <= line + 1;  
        end if;        
      end if;
    end if;
  end process conta_linha;

  -- gera o bitmap
  map1: entity work.ger_palavras port map (key, PS2_DAT, PS2_CLK, CLOCK_24, CLK27M, init_line, init_col, reset, mapaLetras, LEDG, LEDR);
	

  PROCESS (clk27M)
	BEGIN
	
		if reset = '1' then
			pixel_bit <= start_screen(addr);
		elsif clk27M'event and clk27M = '1' then
			IF (col >= init_col AND col < init_col + 5 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 1
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5);
			elsif (col >= init_col + 6 AND col < init_col + 5 + 6 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 2
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 1*(25 - 6));
			elsif (col >= init_col + 12 AND col < init_col + 5 +12 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 3
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 2*(25 - 6));
			elsif (col >= init_col + 18 AND col < init_col + 5 + 18 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 4
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 3*(25 - 6));
			elsif (col >= init_col + 24 AND col < init_col + 29 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 5
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 4*(25 - 6));
			elsif (col >= init_col + 30 AND col < init_col + 35 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 6
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 5*(25 - 6));
			elsif (col >= init_col + 36 AND col < init_col + 41 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 7
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 6*(25 - 6));
			elsif (col >= init_col + 42 AND col < init_col + 47 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 8
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 7*(25 - 6));
			elsif (col >= init_col + 48 AND col < init_col + 53 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 9
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 8*(25 - 6));
			elsif (col >= init_col + 54 AND col < init_col + 59  AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 10 
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 9*(25 - 6));
			elsif (col >= init_col + 60 AND col < init_col + 65 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 11
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 10*(25 - 6));
			elsif (col >= init_col + 66 AND col < init_col + 71 AND line >= init_line AND line < init_line + 5) THEN -- QUADRADO DA LETRA 12
				pixel_bit <= mapaLetras(col - init_col + (line - init_line)*5 + 11*(25 - 6));
			else
				pixel_bit <= '0';
			end if;	
		END IF;	
	END PROCESS;
 
  pixel <= (others => pixel_bit);

  addr  <= col + (128 * line);
  
end comportamento;